magic
tech sky130A
magscale 1 2
timestamp 1605933175
<< nwell >>
rect -382 614 534 910
<< psubdiff >>
rect -150 0 362 96
<< locali >>
rect -153 1291 35 1333
rect -458 1096 -224 1102
rect -458 1016 -320 1096
rect -240 1016 -224 1096
rect -458 1006 -224 1016
rect -458 -49 -408 1006
rect -153 981 -111 1291
rect 322 1167 833 1207
rect -58 1034 -48 1084
rect 2 1034 12 1084
rect -153 939 11 981
rect -31 563 11 939
rect -91 521 33 563
rect -91 442 -49 521
rect 793 447 833 1167
rect -146 400 -49 442
rect 318 428 833 447
rect 314 407 833 428
rect 314 388 376 407
rect -35 -49 15 309
rect -458 -99 15 -49
<< viali >>
rect -320 1016 -240 1096
rect -48 1034 2 1084
<< metal1 >>
rect -610 1384 96 1438
rect -338 1096 -224 1106
rect -338 1016 -320 1096
rect -240 1084 14 1096
rect -240 1034 -48 1084
rect 2 1034 14 1084
rect -240 1016 14 1034
rect -338 1006 -224 1016
rect -610 324 100 378
<< metal2 >>
rect 849 1555 899 1683
rect 693 1505 899 1555
rect 849 98 899 1505
rect 662 92 899 98
rect 588 54 899 92
rect 662 48 899 54
rect 849 -156 899 48
<< metal3 >>
rect 640 684 700 734
rect 706 -156 778 1683
use inverter  inverter_0
timestamp 1604367083
transform 1 0 -332 0 1 446
box -126 -478 242 448
use pass-gate  pass-gate_0
timestamp 1605929851
transform 1 0 210 0 1 218
box -210 -218 503 586
use pass-gate  pass-gate_1
timestamp 1605929851
transform 1 0 210 0 -1 1385
box -210 -218 503 586
<< labels >>
flabel metal1 -588 334 -550 358 0 FreeSans 800 0 0 0 v_in
port 0 nsew
flabel locali 332 396 370 420 0 FreeSans 800 0 0 0 v_out
port 1 nsew
flabel locali -448 110 -410 134 0 FreeSans 800 0 0 0 clk
port 2 nsew
flabel locali -92 408 -54 432 0 FreeSans 800 0 0 0 clk_bar
port 3 nsew
flabel metal3 648 698 686 722 0 FreeSans 800 0 0 0 VPWR
port 4 nsew
flabel metal2 632 58 670 82 0 FreeSans 800 0 0 0 VGND
port 6 nsew
flabel metal1 -592 1392 -560 1420 0 FreeSans 800 0 0 0 v_in2
port 8 nsew
<< end >>
