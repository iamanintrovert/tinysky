* NGSPICE file created from pmos-diff-amp.ext - technology: sky130A

* Include SkyWater sky130 device models
.include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical__lin.spice"
.include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical.spice"
.include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"

* Vdd vdd gnd DC 0.7
* Vgnd vss gnd DC 0.0
* Ibias i_bias vss DC 1n
* Vref in_2 gnd DC 0.3
* Vin in_1 gnd DC 0.2 

Vdd vdd gnd DC 1.8
Vgnd vss gnd DC 0
Ibias i_bias vss DC 1n
Vshort in_2 out DC 0.0
Vin in_1 gnd DC PULSE(0 0.7 100p 0.5u 0.5u 5u 10u)

.subckt sky130_fd_pr__nfet_01v8_r0atdz VSUBS a_n40_n107# a_n98_n81# a_40_n81#
X0 a_40_n81# a_n40_n107# a_n98_n81# VSUBS sky130_fd_pr__nfet_01v8 w=500000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4pknhj VSUBS a_n98_n86# w_n134_n148# a_40_n86# a_n40_n112#
X0 a_40_n86# a_n40_n112# a_n98_n86# w_n134_n148# sky130_fd_pr__pfet_01v8 w=500000u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_4ujh9u VSUBS w_n144_n198# a_n50_n162# a_n108_n136#
+ a_50_n136#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_01v8 w=1e+06u l=500000u
.ends

.subckt pmos-diff-amp in_1 in_2 out i_bias vdd vss
Xsky130_fd_pr__nfet_01v8_r0atdz_0 vss m1_91_n137# m1_91_n137# vss sky130_fd_pr__nfet_01v8_r0atdz
Xsky130_fd_pr__nfet_01v8_r0atdz_1 vss m1_91_n137# vss out sky130_fd_pr__nfet_01v8_r0atdz
Xsky130_fd_pr__pfet_01v8_4pknhj_0 vss m1_91_n137# vdd li_184_186# in_1 sky130_fd_pr__pfet_01v8_4pknhj
Xsky130_fd_pr__pfet_01v8_4ujh9u_0 vss vdd i_bias li_184_186# vdd sky130_fd_pr__pfet_01v8_4ujh9u
Xsky130_fd_pr__pfet_01v8_4pknhj_1 vss li_184_186# vdd out in_2 sky130_fd_pr__pfet_01v8_4pknhj
Xsky130_fd_pr__pfet_01v8_4ujh9u_1 vss vdd i_bias vdd i_bias sky130_fd_pr__pfet_01v8_4ujh9u
.ends

*instantiate
Xdiff in_1 in_2 out i_bias vdd vss pmos-diff-amp

.control
* dc Vin 0 0.7 0.01
* plot v(in_2) v(in_1) v(out)

tran 100n 30u
plot v(in_1) v(out)
.endc
.end


