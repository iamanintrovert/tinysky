* NGSPICE file created from pass-gate-inv.ext - technology: sky130A

* Include SkyWater sky130 device models
.include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical__lin.spice"
.include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical.spice"
.include "/home/mhasan13/pdk/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice"
*.include "/home/mhasan13/pdk/pdk-prepared/sky130A/libs.tech/ngspice/sky130.lib.spice" tt


* DC source for current measure
Vclk clk 0 PULSE(0 1 100p 100p 100p 100n 200n)
Vdd VPWR 0 DC 1.0V
Vgnd VGND 0 DC 0.0V
Vin1 v_in 0 DC 0.2V
Vin2 v_in2 0 DC 0.8V

.subckt sky130_fd_pr__nfet_01v8_8mr83b VSUBS a_n73_n42# a_n15_n68# a_15_n42#
X0 a_15_n42# a_n15_n68# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_ykwexw VSUBS a_n73_n42# w_n109_n104# a_n15_n68# a_15_n42#
X0 a_15_n42# a_n15_n68# a_n73_n42# w_n109_n104# sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends

.subckt inverter GND in VPWR out
Xsky130_fd_pr__nfet_01v8_8mr83b_0 GND GND in out sky130_fd_pr__nfet_01v8_8mr83b
Xsky130_fd_pr__pfet_01v8_ykwexw_0 GND VPWR VPWR in out sky130_fd_pr__pfet_01v8_ykwexw
.ends

.subckt sky130_fd_pr__nfet_01v8_5mkfxl VSUBS a_n73_n42# a_15_n42# a_n33_n130#
X0 a_15_n42# a_n33_n130# a_n73_n42# VSUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_pa2hmj VSUBS a_n33_n177# a_15_n80# w_n109_n180# a_n73_n80#
X0 a_15_n80# a_n33_n177# a_n73_n80# w_n109_n180# sky130_fd_pr__pfet_01v8 w=800000u l=150000u
.ends

.subckt pass-gate clk clk_bar v_in v_out v_newll v_sub
Xsky130_fd_pr__nfet_01v8_5mkfxl_0 v_sub v_out v_in clk sky130_fd_pr__nfet_01v8_5mkfxl
Xsky130_fd_pr__pfet_01v8_pa2hmj_0 v_sub clk_bar v_out v_newll v_in sky130_fd_pr__pfet_01v8_pa2hmj
.ends

.subckt pass-gate-inv v_in v_out clk clk_bar VPWR VGND v_in2
Xinverter_0 VGND clk VPWR clk_bar inverter
Xpass-gate_0 clk clk_bar v_in v_out VPWR VGND pass-gate
Xpass-gate_1 clk_bar clk v_in2 v_out VPWR VGND pass-gate
.ends

Xpass v_in v_out clk clk_bar VPWR VGND v_in2 pass-gate-inv

.control
tran 50p 700n
*dc Vin 0 1 0.01
plot v(clk) v(clk_bar) v(v_out)
.end

.endc

